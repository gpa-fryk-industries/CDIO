library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;


entity audio_mixer is
  generic (
    NUM_CHANNELS: integer := 5;
    CHANNEL_WIDTH: integer := 16
  );
  port (
    -- Basic control
    clk, rst: in std_logic

    --
    




  );
end entity ; -- dds_core

architecture arch_dds_core of dds_core is
  
  
    
begin


end architecture ; -- arch_dds_core


