
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;


package audio_pkg is
	
	subtype s16_audio is signed(15 downto 0);

end package ; -- audio_pkg 





